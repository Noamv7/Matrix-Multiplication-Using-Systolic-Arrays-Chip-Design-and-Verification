`resetall
`timescale 1ns/10ps
